module top();
    input,
    output


    reg;

    
endmodule